module ring_osc(
    output clk_out
);

endmodule