module ring_osc(
    input en,
    
    output clk_out
);

endmodule